module sokol

import shy.wraps.sokol.c as _
import shy.wraps.sokol.f as _
