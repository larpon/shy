module f

import shy.wraps.fontstash
import shy.wraps.sokol.gfx

pub const (
	used_import = fontstash.used_import + gfx.used_import
)
