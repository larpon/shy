// Copyright(C) 2022 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module solid

pub struct Rect {
pub mut:
	x f32
	y f32
	w f32 = 100
	h f32 = 100
}
