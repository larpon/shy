module f

import shy.wraps.fontstash as _
import shy.wraps.sokol.gfx as _
