module sokol

import shy.wraps.sokol.c
import shy.wraps.sokol.f

pub const (
	used_import = c.used_import + f.used_import
)
